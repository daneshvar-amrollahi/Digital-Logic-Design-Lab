library verilog;
use verilog.vl_types.all;
entity ProcessorTB is
end ProcessorTB;
