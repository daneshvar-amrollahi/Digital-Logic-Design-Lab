library verilog;
use verilog.vl_types.all;
entity div113 is
    port(
        output0         : out    vl_logic;
        input3          : in     vl_logic;
        input2          : in     vl_logic;
        input1          : in     vl_logic;
        input0          : in     vl_logic;
        clk             : in     vl_logic;
        preset          : in     vl_logic;
        input7          : in     vl_logic;
        input6          : in     vl_logic;
        input5          : in     vl_logic;
        input4          : in     vl_logic;
        output1         : out    vl_logic;
        output2         : out    vl_logic;
        output3         : out    vl_logic;
        output4         : out    vl_logic;
        output5         : out    vl_logic;
        output6         : out    vl_logic;
        output7         : out    vl_logic;
        MSBcout         : out    vl_logic
    );
end div113;
