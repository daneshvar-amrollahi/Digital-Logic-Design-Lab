library verilog;
use verilog.vl_types.all;
entity WaveGeneratorTB is
end WaveGeneratorTB;
