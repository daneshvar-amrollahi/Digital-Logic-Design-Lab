library verilog;
use verilog.vl_types.all;
entity FreqMult_sv_unit is
end FreqMult_sv_unit;
