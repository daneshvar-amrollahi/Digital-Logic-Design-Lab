library verilog;
use verilog.vl_types.all;
entity count113dispTB is
end count113dispTB;
