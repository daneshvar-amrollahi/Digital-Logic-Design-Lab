library verilog;
use verilog.vl_types.all;
entity CDividerTB is
end CDividerTB;
