library verilog;
use verilog.vl_types.all;
entity exptest is
end exptest;
