library verilog;
use verilog.vl_types.all;
entity FreqMultTB is
end FreqMultTB;
