library verilog;
use verilog.vl_types.all;
entity FuncGenWithFreqSelTB is
end FuncGenWithFreqSelTB;
