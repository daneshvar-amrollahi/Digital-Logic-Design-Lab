library verilog;
use verilog.vl_types.all;
entity FinalTB is
end FinalTB;
