library verilog;
use verilog.vl_types.all;
entity ring_oscill_tb is
end ring_oscill_tb;
