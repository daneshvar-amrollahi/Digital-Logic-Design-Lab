library verilog;
use verilog.vl_types.all;
entity cnt7TB is
end cnt7TB;
