library verilog;
use verilog.vl_types.all;
entity integTB is
end integTB;
