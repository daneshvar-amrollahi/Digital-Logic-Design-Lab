library verilog;
use verilog.vl_types.all;
entity integTB_sv_unit is
end integTB_sv_unit;
