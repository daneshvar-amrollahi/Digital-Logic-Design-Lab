library verilog;
use verilog.vl_types.all;
entity div113tb is
end div113tb;
