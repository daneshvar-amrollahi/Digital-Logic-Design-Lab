library verilog;
use verilog.vl_types.all;
entity lm_555_tb is
end lm_555_tb;
