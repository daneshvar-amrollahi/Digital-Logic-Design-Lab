library verilog;
use verilog.vl_types.all;
entity cnt8TB is
end cnt8TB;
