library verilog;
use verilog.vl_types.all;
entity controller_sv_unit is
end controller_sv_unit;
