library verilog;
use verilog.vl_types.all;
entity integSynTB is
end integSynTB;
