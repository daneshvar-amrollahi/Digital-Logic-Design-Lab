library verilog;
use verilog.vl_types.all;
entity exp2msTB is
end exp2msTB;
